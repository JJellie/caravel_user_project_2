module tb_formal_wishbone (
        input wire clk
);
endmodule